
`timescale 1ns/10ps
parameter GATE_DELAY=0*50.0/1000.0; // 50ns/1000 = 50ps

// Used in testbenches (Adjustable)
parameter TESTBENCH_DELAY=5000;
