
// `define BENCHMARK "benchmarks/test01_AddiB.arm"
// `define BENCHMARK "benchmarks/test02_AddsSubs.arm"
// `define BENCHMARK "benchmarks/test03_CbzB.arm"
// `define BENCHMARK "benchmarks/test04_LdurStur.arm"
// `define BENCHMARK "benchmarks/test05_Blt.arm"
// `define BENCHMARK "benchmarks/test06_MovkMovz.arm"
// `define BENCHMARK "benchmarks/test07_LdurbSturb.arm"
// `define BENCHMARK "benchmarks/test10_forwarding.arm"
// `define BENCHMARK "benchmarks/test11_Sort.arm"
`define BENCHMARK "benchmarks/test12_ToUpper.arm"